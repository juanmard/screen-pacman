// Code for bridge.
module top ( input PIN_22, input CLK,
             output PIN_13, output PIN_12, output PIN_11, output PIN_10, output PIN_9);
    main chimpun (PIN_22, CLK, PIN_13, PIN_12, PIN_11, PIN_10, PIN_9);
endmodule

